`timescale 1ns/10ps

//OOGA BOOGA

module alarm(ss, sp);
    input ss;
    output sp;

    wire ss, sp;
endmodule
